module labM;


